package env_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import my_pkg::*;

  `include "my_env.sv"

endpackage: env_pkg
